module Experimento_2();