module Experimento_1();